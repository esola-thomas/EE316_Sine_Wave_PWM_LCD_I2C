library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity system_state is
port(
	clk : std_logic
	);
end system_state;

architecture arch of system_state is 

begin

end;