entity LCD_Controller is begin

end LCD_Controller;

architecture arch of LCD_Controller is 

begin

end arch;